----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10.01.2018 10:26:09
-- Design Name: 
-- Module Name: RAM2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;



entity RAM2 is

    port (  clk : in std_logic;
    
            adrA : in std_logic_vector (14 - 1 downto 0);
            dOutA : out std_logic_vector (32 - 1 downto 0);
            
            writeEnableB : in std_logic;
            adrB : in std_logic_vector (14 - 1 downto 0);
            dInB : in std_logic_vector (32 - 1 downto 0);
            dOutB : out std_logic_vector (32 - 1 downto 0));

end RAM2;

architecture Behavioral of RAM2 is
type memory_t is array (2**14 - 1 downto 0) of std_logic_vector(32 - 1 downto 0);

constant prog : memory_t :=
(
0=>"00000000000000000001010100010111",
1=>"01001010000001010000010100010011",
2=>"00000000000000001000010110010111",
3=>"11111111100001011000010110010011",
4=>"00000000000000001000011000010111",
5=>"11111111000001100000011000010011",
6=>"00000000000001010010001010000011",
7=>"00000000010001010000010100010011",
8=>"00000000010101011010000000100011",
9=>"00000000010001011000010110010011",
10=>"11111110110001011110100011100011",
11=>"00000000000000001001011000010111",
12=>"11111101010001100000011000010011",
13=>"00000000000001011010000000100011",
14=>"00000000010001011000010110010011",
15=>"11111110101101100111110011100011",
16=>"00000000000000001001000100010111",
17=>"11111100000000010000000100010011",
18=>"00000000000000000000001000010011",
19=>"00000000000000000000000010010011",
20=>"00000000000000000000010000010011",
21=>"01100100110100000000000001101111",
22=>"11111101000000010000000100010011",
23=>"00000010100000010010011000100011",
24=>"00000011000000010000010000010011",
25=>"11111100101001000010111000100011",
26=>"11111100101101000010110000100011",
27=>"00000000000100000000011110010011",
28=>"11111110111101000010011000100011",
29=>"11111110110001000010011100000011",
30=>"11111101100001000010011110000011",
31=>"00000000111101110001011110110011",
32=>"11111110111101000010011000100011",
33=>"11111101110001000010011100000011",
34=>"11111110110001000010011110000011",
35=>"00000000111101110111011110110011",
36=>"00000000000001111001011001100011",
37=>"00000000000000000000011110010011",
38=>"00000000100000000000000001101111",
39=>"00000000000100000000011110010011",
40=>"00000000000001111000010100010011",
41=>"00000010110000010010010000000011",
42=>"00000011000000010000000100010011",
43=>"00000000000000001000000001100111",
44=>"11111101000000010000000100010011",
45=>"00000010100000010010011000100011",
46=>"00000011000000010000010000010011",
47=>"11111100101001000010111000100011",
48=>"11111100101101000010110000100011",
49=>"00000000000100000000011110010011",
50=>"11111110111101000010011000100011",
51=>"11111110110001000010011100000011",
52=>"11111101100001000010011110000011",
53=>"00000000111101110001011110110011",
54=>"11111110111101000010011000100011",
55=>"11111101110001000010011110000011",
56=>"00000000000001111010011100000011",
57=>"11111110110001000010011110000011",
58=>"00000000111101110110011100110011",
59=>"11111101110001000010011110000011",
60=>"00000000111001111010000000100011",
61=>"00000000000000000000000000010011",
62=>"00000010110000010010010000000011",
63=>"00000011000000010000000100010011",
64=>"00000000000000001000000001100111",
65=>"11111101000000010000000100010011",
66=>"00000010100000010010011000100011",
67=>"00000011000000010000010000010011",
68=>"11111100101001000010111000100011",
69=>"11111100101101000010110000100011",
70=>"00000000000100000000011110010011",
71=>"11111110111101000010011000100011",
72=>"11111110110001000010011100000011",
73=>"11111101100001000010011110000011",
74=>"00000000111101110001011110110011",
75=>"11111110111101000010011000100011",
76=>"11111101110001000010011110000011",
77=>"00000000000001111010011100000011",
78=>"11111110110001000010011110000011",
79=>"11111111111101111100011110010011",
80=>"00000000111101110111011100110011",
81=>"11111101110001000010011110000011",
82=>"00000000111001111010000000100011",
83=>"00000000000000000000000000010011",
84=>"00000010110000010010010000000011",
85=>"00000011000000010000000100010011",
86=>"00000000000000001000000001100111",
87=>"11111101000000010000000100010011",
88=>"00000010000100010010011000100011",
89=>"00000010100000010010010000100011",
90=>"00000011000000010000010000010011",
91=>"11111100101001000010111000100011",
92=>"11111100101101000010110000100011",
93=>"11111100110001000010101000100011",
94=>"11111110000001000010011000100011",
95=>"11111101100001000010011110000011",
96=>"11111110111101000010011000100011",
97=>"00000001110000000000000001101111",
98=>"11111110110001000010010110000011",
99=>"11111101110001000010010100000011",
100=>"11110111010111111111000011101111",
101=>"11111110110001000010011110000011",
102=>"00000000000101111000011110010011",
103=>"11111110111101000010011000100011",
104=>"11111110110001000010011100000011",
105=>"11111101010001000010011110000011",
106=>"11111110111001111101000011100011",
107=>"00000000000000000000000000010011",
108=>"00000010110000010010000010000011",
109=>"00000010100000010010010000000011",
110=>"00000011000000010000000100010011",
111=>"00000000000000001000000001100111",
112=>"11111101000000010000000100010011",
113=>"00000010100000010010011000100011",
114=>"00000011000000010000010000010011",
115=>"11111100101001000010111000100011",
116=>"11111100101101000010110000100011",
117=>"11111111111111110000011110110111",
118=>"11111110111101000010011000100011",
119=>"11111110000001000010010000100011",
120=>"11111101110001000010011100000011",
121=>"00000100111100000000011110010011",
122=>"00000000111001111111011001100011",
123=>"00000100111100000000011110010011",
124=>"11111100111101000010111000100011",
125=>"11111101100001000010011100000011",
126=>"00000001110100000000011110010011",
127=>"00000000111001111111011001100011",
128=>"00000001110100000000011110010011",
129=>"11111100111101000010110000100011",
130=>"11111101100001000010011110000011",
131=>"00000000011101111001011110010011",
132=>"11111110111101000010010000100011",
133=>"11111110110001000010011100000011",
134=>"11111110100001000010011110000011",
135=>"00000000111101110000011110110011",
136=>"11111101110001000010011100000011",
137=>"00000000111101110000011110110011",
138=>"11111110111101000010011000100011",
139=>"11111110110001000010011110000011",
140=>"00000000000001111000010100010011",
141=>"00000010110000010010010000000011",
142=>"00000011000000010000000100010011",
143=>"00000000000000001000000001100111",
144=>"11111101000000010000000100010011",
145=>"00000010100000010010011000100011",
146=>"00000011000000010000010000010011",
147=>"11111100101001000010111000100011",
148=>"11111100101101000010110000100011",
149=>"11111110000001000010011000100011",
150=>"11111110000001000010010000100011",
151=>"11111110000001000010010000100011",
152=>"00000010000000000000000001101111",
153=>"11111110110001000010011100000011",
154=>"11111101110001000010011110000011",
155=>"00000000111101110000011110110011",
156=>"11111110111101000010011000100011",
157=>"11111110100001000010011110000011",
158=>"00000000000101111000011110010011",
159=>"11111110111101000010010000100011",
160=>"11111110100001000010011100000011",
161=>"11111101100001000010011110000011",
162=>"11111100111101110100111011100011",
163=>"11111110110001000010011110000011",
164=>"00000000000001111000010100010011",
165=>"00000010110000010010010000000011",
166=>"00000011000000010000000100010011",
167=>"00000000000000001000000001100111",
168=>"11111101000000010000000100010011",
169=>"00000010100000010010011000100011",
170=>"00000011000000010000010000010011",
171=>"11111100101001000010111000100011",
172=>"11111100101101000010110000100011",
173=>"11111100110001000010101000100011",
174=>"11111110000001000010011000100011",
175=>"11111101110001000010011110000011",
176=>"11111110111101000010010000100011",
177=>"11111101100001000010011100000011",
178=>"00000000000100000000011110010011",
179=>"00000110111101110000110001100011",
180=>"11111101100001000010011100000011",
181=>"11111111111100000000011110010011",
182=>"00000110111101110000011001100011",
183=>"11111110100001000010011110000011",
184=>"00000100111100000101100001100011",
185=>"00000010000000000000000001101111",
186=>"11111110110001000010011110000011",
187=>"00000000000101111000011110010011",
188=>"11111110111101000010011000100011",
189=>"11111110100001000010011100000011",
190=>"11111101100001000010011110000011",
191=>"01000000111101110000011110110011",
192=>"11111110111101000010010000100011",
193=>"11111110100001000010011100000011",
194=>"11111101100001000010011110000011",
195=>"11111100111101110101111011100011",
196=>"00000101100000000000000001101111",
197=>"11111110110001000010011110000011",
198=>"00000000000101111000011110010011",
199=>"11111110111101000010011000100011",
200=>"11111110100001000010011100000011",
201=>"11111101100001000010011110000011",
202=>"00000000111101110000011110110011",
203=>"11111110111101000010010000100011",
204=>"11111101100001000010011110000011",
205=>"01000000111100000000011110110011",
206=>"11111110100001000010011100000011",
207=>"11111100111001111101110011100011",
208=>"00000010100000000000000001101111",
209=>"11111101100001000010011100000011",
210=>"00000000000100000000011110010011",
211=>"00000000111101110001100001100011",
212=>"11111110100001000010011110000011",
213=>"11111110111101000010011000100011",
214=>"00000001000000000000000001101111",
215=>"11111110100001000010011110000011",
216=>"01000000111100000000011110110011",
217=>"11111110111101000010011000100011",
218=>"11111101010001000010011110000011",
219=>"00000000000001111000100001100011",
220=>"11111101010001000010011110000011",
221=>"11111110100001000010011100000011",
222=>"00000000111001111010000000100011",
223=>"11111110110001000010011110000011",
224=>"00000000000001111000010100010011",
225=>"00000010110000010010010000000011",
226=>"00000011000000010000000100010011",
227=>"00000000000000001000000001100111",
228=>"11111110000000010000000100010011",
229=>"00000000000100010010111000100011",
230=>"00000000100000010010110000100011",
231=>"00000010000000010000010000010011",
232=>"11111110101001000010011000100011",
233=>"11111110101101000010010000100011",
234=>"11111110110001000010001000100011",
235=>"11111111111111110000011110110111",
236=>"00000001111001111000011110010011",
237=>"11111110111101000010011000100011",
238=>"11111110110001000010011110000011",
239=>"00000010000000000000011100010011",
240=>"00000000111001111010000000100011",
241=>"11111110100001000010011110000011",
242=>"00000100100000000000011100010011",
243=>"00000000111001111010000000100011",
244=>"11111110100001000010011110000011",
245=>"00000110010100000000011100010011",
246=>"00000000111001111010000000100011",
247=>"11111110100001000010011110000011",
248=>"00000111001000000000011100010011",
249=>"00000000111001111010000000100011",
250=>"11111110100001000010011110000011",
251=>"00000111101000000000011100010011",
252=>"00000000111001111010000000100011",
253=>"11111110100001000010011110000011",
254=>"00000110110000000000011100010011",
255=>"00000000111001111010000000100011",
256=>"11111110100001000010011110000011",
257=>"00000110100100000000011100010011",
258=>"00000000111001111010000000100011",
259=>"11111110100001000010011110000011",
260=>"00000110001100000000011100010011",
261=>"00000000111001111010000000100011",
262=>"11111110100001000010011110000011",
263=>"00000110100000000000011100010011",
264=>"00000000111001111010000000100011",
265=>"11111110100001000010011110000011",
266=>"00000000000001111010000000100011",
267=>"11111110100001000010011110000011",
268=>"00000101011100000000011100010011",
269=>"00000000111001111010000000100011",
270=>"11111110100001000010011110000011",
271=>"00000110100100000000011100010011",
272=>"00000000111001111010000000100011",
273=>"11111110100001000010011110000011",
274=>"00000110110000000000011100010011",
275=>"00000000111001111010000000100011",
276=>"11111110100001000010011110000011",
277=>"00000110110000000000011100010011",
278=>"00000000111001111010000000100011",
279=>"11111110100001000010011110000011",
280=>"00000110101100000000011100010011",
281=>"00000000111001111010000000100011",
282=>"11111110100001000010011110000011",
283=>"00000110111100000000011100010011",
284=>"00000000111001111010000000100011",
285=>"11111110100001000010011110000011",
286=>"00000110110100000000011100010011",
287=>"00000000111001111010000000100011",
288=>"11111110100001000010011110000011",
289=>"00000110110100000000011100010011",
290=>"00000000111001111010000000100011",
291=>"11111110100001000010011110000011",
292=>"00000110010100000000011100010011",
293=>"00000000111001111010000000100011",
294=>"11111110100001000010011110000011",
295=>"00000110111000000000011100010011",
296=>"00000000111001111010000000100011",
297=>"11111110100001000010011110000011",
298=>"00000010000100000000011100010011",
299=>"00000000111001111010000000100011",
300=>"11111111111111110000011110110111",
301=>"00011000111101111000011110010011",
302=>"11111110111101000010011000100011",
303=>"11111110110001000010011110000011",
304=>"00000010000000000000011100010011",
305=>"00000000111001111010000000100011",
306=>"11111110100001000010011110000011",
307=>"00000101011100000000011100010011",
308=>"00000000111001111010000000100011",
309=>"11111110100001000010011110000011",
310=>"00000110000100000000011100010011",
311=>"00000000111001111010000000100011",
312=>"11111110100001000010011110000011",
313=>"00000110010100000000011100010011",
314=>"00000000111001111010000000100011",
315=>"11111110100001000010011110000011",
316=>"00000110100000000000011100010011",
317=>"00000000111001111010000000100011",
318=>"11111110100001000010011110000011",
319=>"00000110110000000000011100010011",
320=>"00000000111001111010000000100011",
321=>"11111110100001000010011110000011",
322=>"00000110010100000000011100010011",
323=>"00000000111001111010000000100011",
324=>"11111110100001000010011110000011",
325=>"00000110111000000000011100010011",
326=>"00000000111001111010000000100011",
327=>"11111110100001000010011110000011",
328=>"00000000000001111010000000100011",
329=>"11111110100001000010011110000011",
330=>"00000101001100000000011100010011",
331=>"00000000111001111010000000100011",
332=>"11111110100001000010011110000011",
333=>"00000110100100000000011100010011",
334=>"00000000111001111010000000100011",
335=>"11111110100001000010011110000011",
336=>"00000110010100000000011100010011",
337=>"00000000111001111010000000100011",
338=>"11111110100001000010011110000011",
339=>"00000011101000000000011100010011",
340=>"00000000111001111010000000100011",
341=>"11111111111111110000011110110111",
342=>"00100000111101111000011110010011",
343=>"11111110111101000010011000100011",
344=>"11111110110001000010011110000011",
345=>"00000010000000000000011100010011",
346=>"00000000111001111010000000100011",
347=>"11111110100001000010011110000011",
348=>"00000010110100000000011100010011",
349=>"00000000111001111010000000100011",
350=>"11111110100001000010011110000011",
351=>"00000010000000000000011100010011",
352=>"00000000111001111010000000100011",
353=>"11111110100001000010011110000011",
354=>"00000101001100000000011100010011",
355=>"00000000111001111010000000100011",
356=>"11111110100001000010011110000011",
357=>"00000110100000000000011100010011",
358=>"00000000111001111010000000100011",
359=>"11111110100001000010011110000011",
360=>"00000110111100000000011100010011",
361=>"00000000111001111010000000100011",
362=>"11111110100001000010011110000011",
363=>"00000111011100000000011100010011",
364=>"00000000111001111010000000100011",
365=>"11111111111111110000011110110111",
366=>"00101000111101111000011110010011",
367=>"11111110111101000010011000100011",
368=>"11111110110001000010011110000011",
369=>"00000010000000000000011100010011",
370=>"00000000111001111010000000100011",
371=>"11111110100001000010011110000011",
372=>"00000010110100000000011100010011",
373=>"00000000111001111010000000100011",
374=>"11111110100001000010011110000011",
375=>"00000010000000000000011100010011",
376=>"00000000111001111010000000100011",
377=>"11111110100001000010011110000011",
378=>"00000101010000000000011100010011",
379=>"00000000111001111010000000100011",
380=>"11111110100001000010011110000011",
381=>"00000110000100000000011100010011",
382=>"00000000111001111010000000100011",
383=>"11111110100001000010011110000011",
384=>"00000111001100000000011100010011",
385=>"00000000111001111010000000100011",
386=>"11111110100001000010011110000011",
387=>"00000110001100000000011100010011",
388=>"00000000111001111010000000100011",
389=>"11111110100001000010011110000011",
390=>"00000110100000000000011100010011",
391=>"00000000111001111010000000100011",
392=>"11111110100001000010011110000011",
393=>"00000110010100000000011100010011",
394=>"00000000111001111010000000100011",
395=>"11111110100001000010011110000011",
396=>"00000110111000000000011100010011",
397=>"00000000111001111010000000100011",
398=>"11111110100001000010011110000011",
399=>"00000111001000000000011100010011",
400=>"00000000111001111010000000100011",
401=>"11111110100001000010011110000011",
402=>"00000110010100000000011100010011",
403=>"00000000111001111010000000100011",
404=>"11111110100001000010011110000011",
405=>"00000110001100000000011100010011",
406=>"00000000111001111010000000100011",
407=>"11111110100001000010011110000011",
408=>"00000110100000000000011100010011",
409=>"00000000111001111010000000100011",
410=>"11111110100001000010011110000011",
411=>"00000110111000000000011100010011",
412=>"00000000111001111010000000100011",
413=>"11111110100001000010011110000011",
414=>"00000110010100000000011100010011",
415=>"00000000111001111010000000100011",
416=>"11111110100001000010011110000011",
417=>"00000111001000000000011100010011",
418=>"00000000111001111010000000100011",
419=>"00000001010100000000010110010011",
420=>"00000000011100000000010100010011",
421=>"10110010110111111111000011101111",
422=>"11111110101001000010011000100011",
423=>"11111110110001000010011110000011",
424=>"00000000000001111010000000100011",
425=>"11111110100001000010011110000011",
426=>"00000000011100000000011100010011",
427=>"00000000111001111010000000100011",
428=>"00000001011000000000010110010011",
429=>"00000000010100000000010100010011",
430=>"10110000100111111111000011101111",
431=>"11111110101001000010011000100011",
432=>"11111110110001000010011110000011",
433=>"00000000000001111010000000100011",
434=>"11111110100001000010011110000011",
435=>"00000100100000000000011100010011",
436=>"00000000111001111010000000100011",
437=>"11111110100001000010011110000011",
438=>"00000110111100000000011100010011",
439=>"00000000111001111010000000100011",
440=>"11111110100001000010011110000011",
441=>"00000110001100000000011100010011",
442=>"00000000111001111010000000100011",
443=>"11111110100001000010011110000011",
444=>"00000110100000000000011100010011",
445=>"00000000111001111010000000100011",
446=>"00000001100000000000010110010011",
447=>"00000000001100000000010100010011",
448=>"10101100000111111111000011101111",
449=>"11111110101001000010011000100011",
450=>"11111110110001000010011110000011",
451=>"00000000000001111010000000100011",
452=>"11111110100001000010011110000011",
453=>"00000000011100000000011100010011",
454=>"00000000111001111010000000100011",
455=>"11111110100001000010011110000011",
456=>"00000000000001111010000000100011",
457=>"11111110100001000010011110000011",
458=>"00000000000001111010000000100011",
459=>"11111110100001000010011110000011",
460=>"00000000000001111010000000100011",
461=>"11111110100001000010011110000011",
462=>"00000000011100000000011100010011",
463=>"00000000111001111010000000100011",
464=>"11111110100001000010011110000011",
465=>"00000000000001111010000000100011",
466=>"11111110100001000010011110000011",
467=>"00000000000001111010000000100011",
468=>"11111110100001000010011110000011",
469=>"00000000000001111010000000100011",
470=>"11111110100001000010011110000011",
471=>"00000000011100000000011100010011",
472=>"00000000111001111010000000100011",
473=>"00000001100100000000010110010011",
474=>"00000000010100000000010100010011",
475=>"10100101010111111111000011101111",
476=>"11111110101001000010011000100011",
477=>"11111110110001000010011110000011",
478=>"00000000000001111010000000100011",
479=>"11111110100001000010011110000011",
480=>"00000100010100000000011100010011",
481=>"00000000111001111010000000100011",
482=>"11111110100001000010011110000011",
483=>"00000110111000000000011100010011",
484=>"00000000111001111010000000100011",
485=>"11111110100001000010011110000011",
486=>"00000111010000000000011100010011",
487=>"00000000111001111010000000100011",
488=>"11111110100001000010011110000011",
489=>"00000110010100000000011100010011",
490=>"00000000111001111010000000100011",
491=>"11111110100001000010011110000011",
492=>"00000111001000000000011100010011",
493=>"00000000111001111010000000100011",
494=>"00000001101100000000010110010011",
495=>"00000000011100000000010100010011",
496=>"10100000000111111111000011101111",
497=>"11111110101001000010011000100011",
498=>"11111110110001000010011110000011",
499=>"00000000000001111010000000100011",
500=>"11111110100001000010011110000011",
501=>"00000000011100000000011100010011",
502=>"00000000111001111010000000100011",
503=>"00000001110000000000010110010011",
504=>"00000000010100000000010100010011",
505=>"10011101110111111111000011101111",
506=>"11111110101001000010011000100011",
507=>"11111110110001000010011110000011",
508=>"00000000000001111010000000100011",
509=>"11111110100001000010011110000011",
510=>"00000101001000000000011100010011",
511=>"00000000111001111010000000100011",
512=>"11111110100001000010011110000011",
513=>"00000111010100000000011100010011",
514=>"00000000111001111010000000100011",
515=>"11111110100001000010011110000011",
516=>"00000110111000000000011100010011",
517=>"00000000111001111010000000100011",
518=>"11111110100001000010011110000011",
519=>"00000111010000000000011100010011",
520=>"00000000111001111010000000100011",
521=>"11111110100001000010011110000011",
522=>"00000110010100000000011100010011",
523=>"00000000111001111010000000100011",
524=>"11111110100001000010011110000011",
525=>"00000111001000000000011100010011",
526=>"00000000111001111010000000100011",
527=>"00000000010000000000010110010011",
528=>"00000000111100000000010100010011",
529=>"10010111110111111111000011101111",
530=>"11111110101001000010011000100011",
531=>"00000000000000000000000000010011",
532=>"00000001110000010010000010000011",
533=>"00000001100000010010010000000011",
534=>"00000010000000010000000100010011",
535=>"00000000000000001000000001100111",
536=>"11111101000000010000000100010011",
537=>"00000010100000010010011000100011",
538=>"00000011000000010000010000010011",
539=>"11111100101001000010111000100011",
540=>"11111100101101000010110000100011",
541=>"11111100110001000010101000100011",
542=>"11111101110001000010011110000011",
543=>"00000000000001111010000000100011",
544=>"11111110000001000010011000100011",
545=>"00000100000000000000000001101111",
546=>"11111110000001000010010000100011",
547=>"00000001100000000000000001101111",
548=>"11111101100001000010011110000011",
549=>"00000000000001111010000000100011",
550=>"11111110100001000010011110000011",
551=>"00000000000101111000011110010011",
552=>"11111110111101000010010000100011",
553=>"11111110100001000010011100000011",
554=>"00000100111100000000011110010011",
555=>"11111110111001111101001011100011",
556=>"11111101010001000010011110000011",
557=>"00000000000001111010000000100011",
558=>"11111110110001000010011110000011",
559=>"00000000000101111000011110010011",
560=>"11111110111101000010011000100011",
561=>"11111110110001000010011100000011",
562=>"00000001110100000000011110010011",
563=>"11111010111001111101111011100011",
564=>"00000000000000000000000000010011",
565=>"00000010110000010010010000000011",
566=>"00000011000000010000000100010011",
567=>"00000000000000001000000001100111",
568=>"11111110000000010000000100010011",
569=>"00000000000100010010111000100011",
570=>"00000000100000010010110000100011",
571=>"00000010000000010000010000010011",
572=>"11111110101001000010011000100011",
573=>"11111110101101000010010000100011",
574=>"00000000000000000000000000010011",
575=>"11111110100001000010011110000011",
576=>"00000000000001111010011110000011",
577=>"11111110110001000010010110000011",
578=>"00000000000001111000010100010011",
579=>"11110100110011111111000011101111",
580=>"00000000000001010000011100010011",
581=>"00000000000100000000011110010011",
582=>"11111110111101110000001011100011",
583=>"00000000000000000000000000010011",
584=>"00000001110000010010000010000011",
585=>"00000001100000010010010000000011",
586=>"00000010000000010000000100010011",
587=>"00000000000000001000000001100111",
588=>"11111110000000010000000100010011",
589=>"00000000000100010010111000100011",
590=>"00000000100000010010110000100011",
591=>"00000010000000010000010000010011",
592=>"11111110101001000010011000100011",
593=>"11111110101101000010010000100011",
594=>"11111110110001000010001000100011",
595=>"00000000111000000000010110010011",
596=>"00000010000100000000010100010011",
597=>"10000110110111111111000011101111",
598=>"11111110101001000010011000100011",
599=>"11111110110001000010011110000011",
600=>"00000000000001111010000000100011",
601=>"11111110100001000010011110000011",
602=>"00000100100000000000011100010011",
603=>"00000000111001111010000000100011",
604=>"11111110100001000010011110000011",
605=>"00000110010100000000011100010011",
606=>"00000000111001111010000000100011",
607=>"11111110100001000010011110000011",
608=>"00000110110000000000011100010011",
609=>"00000000111001111010000000100011",
610=>"11111110100001000010011110000011",
611=>"00000110110000000000011100010011",
612=>"00000000111001111010000000100011",
613=>"11111110100001000010011110000011",
614=>"00000110111100000000011100010011",
615=>"00000000111001111010000000100011",
616=>"11111110100001000010011110000011",
617=>"00000010000000000000011100010011",
618=>"00000000111001111010000000100011",
619=>"11111110100001000010011110000011",
620=>"00000101011100000000011100010011",
621=>"00000000111001111010000000100011",
622=>"11111110100001000010011110000011",
623=>"00000110111100000000011100010011",
624=>"00000000111001111010000000100011",
625=>"11111110100001000010011110000011",
626=>"00000111001000000000011100010011",
627=>"00000000111001111010000000100011",
628=>"11111110100001000010011110000011",
629=>"00000110110000000000011100010011",
630=>"00000000111001111010000000100011",
631=>"11111110100001000010011110000011",
632=>"00000110010000000000011100010011",
633=>"00000000111001111010000000100011",
634=>"11111110100001000010011110000011",
635=>"00000010000100000000011100010011",
636=>"00000000111001111010000000100011",
637=>"11111110100001000010011110000011",
638=>"00000000001100000000011100010011",
639=>"00000000111001111010000000100011",
640=>"00000001010100000000010110010011",
641=>"00000000011100000000010100010011",
642=>"11111011100011111111000011101111",
643=>"11111110101001000010011000100011",
644=>"11111110110001000010011110000011",
645=>"00000000000001111010000000100011",
646=>"11111110100001000010011110000011",
647=>"00000000011100000000011100010011",
648=>"00000000111001111010000000100011",
649=>"00000001100000000000010110010011",
650=>"00000000001100000000010100010011",
651=>"11111001010011111111000011101111",
652=>"11111110101001000010011000100011",
653=>"11111110110001000010011110000011",
654=>"00000000000001111010000000100011",
655=>"11111110100001000010011110000011",
656=>"00000000011100000000011100010011",
657=>"00000000111001111010000000100011",
658=>"11111110100001000010011110000011",
659=>"00000000000001111010000000100011",
660=>"11111110100001000010011110000011",
661=>"00000000000001111010000000100011",
662=>"11111110100001000010011110000011",
663=>"00000000000001111010000000100011",
664=>"11111110100001000010011110000011",
665=>"00000000011100000000011100010011",
666=>"00000000111001111010000000100011",
667=>"11111110100001000010011110000011",
668=>"00000000000001111010000000100011",
669=>"11111110100001000010011110000011",
670=>"00000000000001111010000000100011",
671=>"11111110100001000010011110000011",
672=>"00000000000001111010000000100011",
673=>"11111110100001000010011110000011",
674=>"00000000011100000000011100010011",
675=>"00000000111001111010000000100011",
676=>"00000001100100000000010110010011",
677=>"00000000010100000000010100010011",
678=>"11110010100011111111000011101111",
679=>"11111110101001000010011000100011",
680=>"11111110110001000010011110000011",
681=>"00000000000001111010000000100011",
682=>"11111110100001000010011110000011",
683=>"00000100001000000000011100010011",
684=>"00000000111001111010000000100011",
685=>"11111110100001000010011110000011",
686=>"00000110000100000000011100010011",
687=>"00000000111001111010000000100011",
688=>"11111110100001000010011110000011",
689=>"00000110001100000000011100010011",
690=>"00000000111001111010000000100011",
691=>"11111110100001000010011110000011",
692=>"00000110101100000000011100010011",
693=>"00000000111001111010000000100011",
694=>"00000001101100000000010110010011",
695=>"00000000011100000000010100010011",
696=>"11101110000011111111000011101111",
697=>"11111110101001000010011000100011",
698=>"11111110110001000010011110000011",
699=>"00000000000001111010000000100011",
700=>"11111110100001000010011110000011",
701=>"00000000011100000000011100010011",
702=>"00000000111001111010000000100011",
703=>"00000000000000000000000000010011",
704=>"00000001110000010010000010000011",
705=>"00000001100000010010010000000011",
706=>"00000010000000010000000100010011",
707=>"00000000000000001000000001100111",
708=>"11111110000000010000000100010011",
709=>"00000000000100010010111000100011",
710=>"00000000100000010010110000100011",
711=>"00000010000000010000010000010011",
712=>"11111110101001000010011000100011",
713=>"11111110101101000010010000100011",
714=>"11111110110001000010001000100011",
715=>"00000000000000000000010110010011",
716=>"00000010000100000000010100010011",
717=>"11101000110011111111000011101111",
718=>"11111110101001000010011000100011",
719=>"11111110110001000010011110000011",
720=>"00000000000001111010000000100011",
721=>"11111110100001000010011110000011",
722=>"00000101010000000000011100010011",
723=>"00000000111001111010000000100011",
724=>"11111110100001000010011110000011",
725=>"00000110000100000000011100010011",
726=>"00000000111001111010000000100011",
727=>"11111110100001000010011110000011",
728=>"00000111001100000000011100010011",
729=>"00000000111001111010000000100011",
730=>"11111110100001000010011110000011",
731=>"00000110001100000000011100010011",
732=>"00000000111001111010000000100011",
733=>"11111110100001000010011110000011",
734=>"00000110100000000000011100010011",
735=>"00000000111001111010000000100011",
736=>"11111110100001000010011110000011",
737=>"00000110010100000000011100010011",
738=>"00000000111001111010000000100011",
739=>"11111110100001000010011110000011",
740=>"00000110111000000000011100010011",
741=>"00000000111001111010000000100011",
742=>"11111110100001000010011110000011",
743=>"00000111001000000000011100010011",
744=>"00000000111001111010000000100011",
745=>"11111110100001000010011110000011",
746=>"00000110010100000000011100010011",
747=>"00000000111001111010000000100011",
748=>"11111110100001000010011110000011",
749=>"00000110001100000000011100010011",
750=>"00000000111001111010000000100011",
751=>"11111110100001000010011110000011",
752=>"00000110100000000000011100010011",
753=>"00000000111001111010000000100011",
754=>"11111110100001000010011110000011",
755=>"00000110111000000000011100010011",
756=>"00000000111001111010000000100011",
757=>"11111110100001000010011110000011",
758=>"00000110010100000000011100010011",
759=>"00000000111001111010000000100011",
760=>"11111110100001000010011110000011",
761=>"00000111001000000000011100010011",
762=>"00000000111001111010000000100011",
763=>"00000001010100000000010110010011",
764=>"00000000011100000000010100010011",
765=>"11011100110011111111000011101111",
766=>"11111110101001000010011000100011",
767=>"11111110110001000010011110000011",
768=>"00000000000001111010000000100011",
769=>"11111110100001000010011110000011",
770=>"00000000011100000000011100010011",
771=>"00000000111001111010000000100011",
772=>"00000001100000000000010110010011",
773=>"00000000001100000000010100010011",
774=>"11011010100011111111000011101111",
775=>"11111110101001000010011000100011",
776=>"11111110110001000010011110000011",
777=>"00000000000001111010000000100011",
778=>"11111110100001000010011110000011",
779=>"00000000011100000000011100010011",
780=>"00000000111001111010000000100011",
781=>"11111110100001000010011110000011",
782=>"00000000000001111010000000100011",
783=>"11111110100001000010011110000011",
784=>"00000000000001111010000000100011",
785=>"11111110100001000010011110000011",
786=>"00000000000001111010000000100011",
787=>"11111110100001000010011110000011",
788=>"00000000011100000000011100010011",
789=>"00000000111001111010000000100011",
790=>"11111110100001000010011110000011",
791=>"00000000000001111010000000100011",
792=>"11111110100001000010011110000011",
793=>"00000000000001111010000000100011",
794=>"11111110100001000010011110000011",
795=>"00000000000001111010000000100011",
796=>"11111110100001000010011110000011",
797=>"00000000011100000000011100010011",
798=>"00000000111001111010000000100011",
799=>"00000001100100000000010110010011",
800=>"00000000000100000000010100010011",
801=>"11010011110011111111000011101111",
802=>"11111110101001000010011000100011",
803=>"11111110110001000010011110000011",
804=>"00000000000001111010000000100011",
805=>"11111110100001000010011110000011",
806=>"00000100001000000000011100010011",
807=>"00000000111001111010000000100011",
808=>"11111110100001000010011110000011",
809=>"00000110000100000000011100010011",
810=>"00000000111001111010000000100011",
811=>"11111110100001000010011110000011",
812=>"00000110001100000000011100010011",
813=>"00000000111001111010000000100011",
814=>"11111110100001000010011110000011",
815=>"00000110101100000000011100010011",
816=>"00000000111001111010000000100011",
817=>"11111110100001000010011110000011",
818=>"00000000000001111010000000100011",
819=>"11111110100001000010011110000011",
820=>"00000000000001111010000000100011",
821=>"11111110100001000010011110000011",
822=>"00000000000001111010000000100011",
823=>"11111110100001000010011110000011",
824=>"00000000000001111010000000100011",
825=>"11111110100001000010011110000011",
826=>"00000000000001111010000000100011",
827=>"11111110100001000010011110000011",
828=>"00000100010100000000011100010011",
829=>"00000000111001111010000000100011",
830=>"11111110100001000010011110000011",
831=>"00000110111000000000011100010011",
832=>"00000000111001111010000000100011",
833=>"11111110100001000010011110000011",
834=>"00000111010000000000011100010011",
835=>"00000000111001111010000000100011",
836=>"11111110100001000010011110000011",
837=>"00000110010100000000011100010011",
838=>"00000000111001111010000000100011",
839=>"11111110100001000010011110000011",
840=>"00000111001000000000011100010011",
841=>"00000000111001111010000000100011",
842=>"00000001101100000000010110010011",
843=>"00000000011100000000010100010011",
844=>"11001001000011111111000011101111",
845=>"11111110101001000010011000100011",
846=>"11111110110001000010011110000011",
847=>"00000000000001111010000000100011",
848=>"11111110100001000010011110000011",
849=>"00000000011100000000011100010011",
850=>"00000000111001111010000000100011",
851=>"00000000000000000000000000010011",
852=>"00000001110000010010000010000011",
853=>"00000001100000010010010000000011",
854=>"00000010000000010000000100010011",
855=>"00000000000000001000000001100111",
856=>"11111010000000010000000100010011",
857=>"00000100000100010010111000100011",
858=>"00000100100000010010110000100011",
859=>"00000110000000010000010000010011",
860=>"11111010101001000010011000100011",
861=>"11111010101101000010010000100011",
862=>"11111010110001000010011110000011",
863=>"11111110111101000010000000100011",
864=>"11111110000001000010001000100011",
865=>"00111011100110101101011110110111",
866=>"10100000000001111000011110010011",
867=>"11111010111101000010110000100011",
868=>"00000101111101011110011110110111",
869=>"00010000000001111000011110010011",
870=>"11111010111101000010111000100011",
871=>"00000000100110001001011110110111",
872=>"01101000000001111000011110010011",
873=>"11111100111101000010000000100011",
874=>"00000000000011110100011110110111",
875=>"00100100000001111000011110010011",
876=>"11111100111101000010001000100011",
877=>"00000000000000011000011110110111",
878=>"01101010000001111000011110010011",
879=>"11111100111101000010010000100011",
880=>"00000000000000000010011110110111",
881=>"01110001000001111000011110010011",
882=>"11111100111101000010011000100011",
883=>"00111110100000000000011110010011",
884=>"11111100111101000010100000100011",
885=>"00000110010000000000011110010011",
886=>"11111100111101000010101000100011",
887=>"00000000101000000000011110010011",
888=>"11111100111101000010110000100011",
889=>"00000000000100000000011110010011",
890=>"11111100111101000010111000100011",
891=>"11111110000001000010010000100011",
892=>"11111010110001000010011110000011",
893=>"00000000000001111101100001100011",
894=>"11111010100001000010011110000011",
895=>"00000010110100000000011100010011",
896=>"00000000111001111010000000100011",
897=>"11111110000001000010011000100011",
898=>"00000111100000000000000001101111",
899=>"11111110000001000010011100000011",
900=>"11111110110001000010011110000011",
901=>"00000000001001111001011110010011",
902=>"11111111000001000000011010010011",
903=>"00000000111101101000011110110011",
904=>"11111100100001111010011110000011",
905=>"11111110000001000000011010010011",
906=>"00000000000001101000011000010011",
907=>"00000000000001111000010110010011",
908=>"00000000000001110000010100010011",
909=>"11000110110011111111000011101111",
910=>"11111110101001000010001000100011",
911=>"11111110100001000010011110000011",
912=>"00000000000001111001110001100011",
913=>"11111110010001000010011110000011",
914=>"00000000000001111001100001100011",
915=>"11111110110001000010011100000011",
916=>"00000000100100000000011110010011",
917=>"00000010111101110001000001100011",
918=>"11111110010001000010011110000011",
919=>"00000011000001111000011110010011",
920=>"00000000000001111000011100010011",
921=>"11111010100001000010011110000011",
922=>"00000000111001111010000000100011",
923=>"00000000000100000000011110010011",
924=>"11111110111101000010010000100011",
925=>"11111110110001000010011110000011",
926=>"00000000000101111000011110010011",
927=>"11111110111101000010011000100011",
928=>"11111110110001000010011100000011",
929=>"00000000100100000000011110010011",
930=>"11111000111001111101001011100011",
931=>"00000000000000000000000000010011",
932=>"00000101110000010010000010000011",
933=>"00000101100000010010010000000011",
934=>"00000110000000010000000100010011",
935=>"00000000000000001000000001100111",
936=>"11111011000000010000000100010011",
937=>"00000100000100010010011000100011",
938=>"00000100100000010010010000100011",
939=>"00000101000000010000010000010011",
940=>"11111111111111111000011110110111",
941=>"11111100111101000010100000100011",
942=>"11111111111111111100011110110111",
943=>"11111100111101000010011000100011",
944=>"11111111111111110000011110110111",
945=>"11111100111101000010010000100011",
946=>"11111111111111110000011110110111",
947=>"11111110111101000010011000100011",
948=>"10000000000000000000011110110111",
949=>"11111100111101000010001000100011",
950=>"10000000000000000000011110110111",
951=>"00000000000101111000011110010011",
952=>"11111100111101000010000000100011",
953=>"11111110000001000010010000100011",
954=>"00000000000100000000011110010011",
955=>"11111110111101000010001000100011",
956=>"11111010000001000010110000100011",
957=>"11111110000001000010000000100011",
958=>"11111100000001000010111000100011",
959=>"11111010000001000010101000100011",
960=>"11111010000001000010111000100011",
961=>"11111100000001000010110000100011",
962=>"11111100000001000010101000100011",
963=>"11111100000001000010011110000011",
964=>"00000000000001111010011100000011",
965=>"11111100010001000010011110000011",
966=>"00000000111001111010000000100011",
967=>"11111101000001000010011110000011",
968=>"00000110010100000000011100010011",
969=>"00000000111001111010000000100011",
970=>"11111110100001000010011110000011",
971=>"00000000000100000000011100010011",
972=>"00010100111001111000100001100011",
973=>"00000000001000000000011100010011",
974=>"00011010111001111000111001100011",
975=>"01010100000001111001000001100011",
976=>"11111110010001000010011110000011",
977=>"00000010000001111000010001100011",
978=>"11111100110001000010011000000011",
979=>"11111101000001000010010110000011",
980=>"11111100100001000010010100000011",
981=>"10010000110111111111000011101111",
982=>"11111100110001000010011000000011",
983=>"11111101000001000010010110000011",
984=>"11111110110001000010010100000011",
985=>"11000010110011111111000011101111",
986=>"11111110000001000010001000100011",
987=>"11111100000001000010011110000011",
988=>"00000000000001111010011110000011",
989=>"11111010111101000010110000100011",
990=>"11111011100001000010011110000011",
991=>"00000001000000000000010110010011",
992=>"00000000000001111000010100010011",
993=>"10001101010011111111000011101111",
994=>"00000000000001010000011100010011",
995=>"00000000000100000000011110010011",
996=>"00000000111101110001111001100011",
997=>"11111110000001000010011110000011",
998=>"00000000000101111000011110010011",
999=>"11111110111101000010010000100011",
1000=>"11111100000001000010010110000011",
1001=>"00000001000000000000010100010011",
1002=>"10010011100111111111000011101111",
1003=>"11111011100001000010011110000011",
1004=>"00000001000100000000010110010011",
1005=>"00000000000001111000010100010011",
1006=>"10001010000011111111000011101111",
1007=>"00000000000001010000011100010011",
1008=>"00000000000100000000011110010011",
1009=>"00000100111101110001100001100011",
1010=>"11111110000001000010011110000011",
1011=>"11111111111101111000011110010011",
1012=>"11111110111101000010000000100011",
1013=>"11111100000001000010010110000011",
1014=>"00000001000100000000010100010011",
1015=>"10010000010111111111000011101111",
1016=>"11111110000001000010011110000011",
1017=>"00000010000001111101000001100011",
1018=>"00000000000100000000011110010011",
1019=>"11111110111101000010000000100011",
1020=>"00000000010100000000010110010011",
1021=>"00000000111100000000010100010011",
1022=>"10011100100011111111000011101111",
1023=>"11111110101001000010011000100011",
1024=>"00000001010000000000000001101111",
1025=>"00000000010000000000010110010011",
1026=>"00000000111100000000010100010011",
1027=>"10011011010011111111000011101111",
1028=>"11111110101001000010011000100011",
1029=>"11111011100001000010011110000011",
1030=>"00000001001000000000010110010011",
1031=>"00000000000001111000010100010011",
1032=>"10000011100011111111000011101111",
1033=>"00000000000001010000011100010011",
1034=>"00000000000100000000011110010011",
1035=>"01000100111101110001110001100011",
1036=>"11111110000001000010011110000011",
1037=>"00000000000101111000011110010011",
1038=>"11111110111101000010000000100011",
1039=>"11111100000001000010010110000011",
1040=>"00000001001000000000010100010011",
1041=>"10001001110111111111000011101111",
1042=>"11111110000001000010011100000011",
1043=>"00000000000100000000011110010011",
1044=>"00000000111001111101111001100011",
1045=>"11111110000001000010000000100011",
1046=>"00000000010000000000010110010011",
1047=>"00000000111100000000010100010011",
1048=>"10010110000011111111000011101111",
1049=>"11111110101001000010011000100011",
1050=>"01000001110000000000000001101111",
1051=>"00000000010100000000010110010011",
1052=>"00000000111100000000010100010011",
1053=>"10010100110011111111000011101111",
1054=>"11111110101001000010011000100011",
1055=>"01000000100000000000000001101111",
1056=>"11111110010001000010011100000011",
1057=>"00000000000100000000011110010011",
1058=>"00000010111101110000011001100011",
1059=>"11111100110001000010011000000011",
1060=>"11111101000001000010010110000011",
1061=>"11111100100001000010010100000011",
1062=>"11111100100011111111000011101111",
1063=>"11111100110001000010011000000011",
1064=>"11111101000001000010010110000011",
1065=>"11111110110001000010010100000011",
1066=>"10001000100111111111000011101111",
1067=>"00000000000100000000011110010011",
1068=>"11111110111101000010001000100011",
1069=>"11111100000001000010011110000011",
1070=>"00000000000001111010011110000011",
1071=>"11111010111101000010110000100011",
1072=>"11111011100001000010011110000011",
1073=>"00000001000000000000010110010011",
1074=>"00000000000001111000010100010011",
1075=>"11111000110111111110000011101111",
1076=>"00000000000001010000011100010011",
1077=>"00000000000100000000011110010011",
1078=>"00111010111101110001101001100011",
1079=>"11111110000001000010010000100011",
1080=>"11111100000001000010010110000011",
1081=>"00000001000000000000010100010011",
1082=>"11111111100011111111000011101111",
1083=>"11111110000001000010000000100011",
1084=>"00111001110000000000000001101111",
1085=>"11111110010001000010011100000011",
1086=>"00000000001000000000011110010011",
1087=>"00000010111101110000011001100011",
1088=>"11111100110001000010011000000011",
1089=>"11111101000001000010010110000011",
1090=>"11111100100001000010010100000011",
1091=>"11110101010011111111000011101111",
1092=>"11111100110001000010011000000011",
1093=>"11111101000001000010010110000011",
1094=>"11111110110001000010010100000011",
1095=>"10011111010111111111000011101111",
1096=>"00000000001000000000011110010011",
1097=>"11111110111101000010001000100011",
1098=>"11111100000001000010011110000011",
1099=>"00000000000001111010011110000011",
1100=>"11111010111101000010110000100011",
1101=>"11111011100001000010011110000011",
1102=>"00000001001100000000010110010011",
1103=>"00000000000001111000010100010011",
1104=>"11110001100111111110000011101111",
1105=>"00000000000001010000011100010011",
1106=>"00000000000100000000011110010011",
1107=>"00000000111101110001111001100011",
1108=>"11111110000001000010010000100011",
1109=>"11111100000001000010010110000011",
1110=>"00000001001100000000010100010011",
1111=>"11111000010011111111000011101111",
1112=>"11111110000001000010000000100011",
1113=>"11111100000001000010111000100011",
1114=>"11111011100001000010011110000011",
1115=>"00000001010000000000010110010011",
1116=>"00000000000001111000010100010011",
1117=>"11101110010111111110000011101111",
1118=>"00000000000001010000011100010011",
1119=>"00000000000100000000011110010011",
1120=>"11011010111101110001010011100011",
1121=>"11111100000001000010010110000011",
1122=>"00000001010000000000010100010011",
1123=>"11110101010011111111000011101111",
1124=>"11111100000001000010011110000011",
1125=>"00000000000001111010011100000011",
1126=>"11111100010001000010011110000011",
1127=>"00000000111001111010000000100011",
1128=>"11111101110001000010011110000011",
1129=>"00000000000100000000011100010011",
1130=>"00000110111001111000011001100011",
1131=>"00000000001000000000011100010011",
1132=>"00010000111001111000110001100011",
1133=>"00101000000001111001111001100011",
1134=>"11111011100001000000011110010011",
1135=>"00000001010000000000010110010011",
1136=>"00000000000001111000010100010011",
1137=>"11110100000111111110000011101111",
1138=>"11111100000001000010011110000011",
1139=>"00000000000001111010011110000011",
1140=>"11111010111101000010101000100011",
1141=>"11111101110001000010011110000011",
1142=>"00000000000101111000011110010011",
1143=>"11111100111101000010111000100011",
1144=>"00000000010100000000010110010011",
1145=>"00000001010000000000010100010011",
1146=>"11111101100111111110000011101111",
1147=>"11111110101001000010011000100011",
1148=>"11111110110001000010011110000011",
1149=>"00000000000001111010000000100011",
1150=>"11111011010001000010011110000011",
1151=>"11111101000001000010010110000011",
1152=>"00000000000001111000010100010011",
1153=>"10110101110111111111000011101111",
1154=>"11111101000001000010011110000011",
1155=>"00000000000001111010000000100011",
1156=>"00100110100000000000000001101111",
1157=>"11111011100001000000011110010011",
1158=>"00000001010000000000010110010011",
1159=>"00000000000001111000010100010011",
1160=>"11101110010111111110000011101111",
1161=>"11111100000001000010011110000011",
1162=>"00000000000001111010011110000011",
1163=>"11111100111101000010110000100011",
1164=>"11111101110001000010011110000011",
1165=>"00000000000101111000011110010011",
1166=>"11111100111101000010111000100011",
1167=>"11111101100001000010011110000011",
1168=>"00000000000100000000011100010011",
1169=>"00000010111001111000110001100011",
1170=>"00000000000100000000011100010011",
1171=>"00000000111101110100011001100011",
1172=>"00000000000001111000111001100011",
1173=>"00000101100000000000000001101111",
1174=>"00000000001000000000011100010011",
1175=>"00000010111001111000100001100011",
1176=>"00000000001100000000011100010011",
1177=>"00000010111001111000110001100011",
1178=>"00000100010000000000000001101111",
1179=>"11111101000001000010011110000011",
1180=>"00000010101100000000011100010011",
1181=>"00000000111001111010000000100011",
1182=>"00000100010000000000000001101111",
1183=>"11111101000001000010011110000011",
1184=>"00000010110100000000011100010011",
1185=>"00000000111001111010000000100011",
1186=>"00000011010000000000000001101111",
1187=>"11111101000001000010011110000011",
1188=>"00000010101000000000011100010011",
1189=>"00000000111001111010000000100011",
1190=>"00000010010000000000000001101111",
1191=>"11111101000001000010011110000011",
1192=>"00000010111100000000011100010011",
1193=>"00000000111001111010000000100011",
1194=>"00000001010000000000000001101111",
1195=>"11111101000001000010011110000011",
1196=>"00000010010100000000011100010011",
1197=>"00000000111001111010000000100011",
1198=>"00000000000000000000000000010011",
1199=>"11111101000001000010011110000011",
1200=>"00000000000001111010000000100011",
1201=>"00011011010000000000000001101111",
1202=>"11111011100001000000011110010011",
1203=>"00000001111100000000011000010011",
1204=>"00000001000000000000010110010011",
1205=>"00000000000001111000010100010011",
1206=>"11101000010111111110000011101111",
1207=>"11111100000001000010011110000011",
1208=>"00000000000001111010011110000011",
1209=>"11111010111101000010111000100011",
1210=>"11111101110001000010011110000011",
1211=>"00000000000101111000011110010011",
1212=>"11111100111101000010111000100011",
1213=>"11111101000001000010010110000011",
1214=>"11111011110001000010010100000011",
1215=>"10100110010111111111000011101111",
1216=>"11111101000001000010011110000011",
1217=>"00000000000001111010000000100011",
1218=>"11111101000001000010011110000011",
1219=>"00000011110100000000011100010011",
1220=>"00000000111001111010000000100011",
1221=>"11111101000001000010011110000011",
1222=>"00000000000001111010000000100011",
1223=>"11111101100001000010011110000011",
1224=>"00000000000100000000011100010011",
1225=>"00000010111001111000111001100011",
1226=>"00000000000100000000011100010011",
1227=>"00000000111101110100011001100011",
1228=>"00000000000001111000111001100011",
1229=>"00001001000000000000000001101111",
1230=>"00000000001000000000011100010011",
1231=>"00000010111001111000110001100011",
1232=>"00000000001100000000011100010011",
1233=>"00000100111001111000011001100011",
1234=>"00000111110000000000000001101111",
1235=>"11111011010001000010011100000011",
1236=>"11111011110001000010011110000011",
1237=>"00000000111101110000011110110011",
1238=>"11111010111101000010101000100011",
1239=>"00001001100000000000000001101111",
1240=>"11111011010001000010011100000011",
1241=>"11111011110001000010011110000011",
1242=>"01000000111101110000011110110011",
1243=>"11111010111101000010101000100011",
1244=>"00001000010000000000000001101111",
1245=>"11111011010001000010011110000011",
1246=>"11111011110001000010010110000011",
1247=>"00000000000001111000010100010011",
1248=>"11101100000111111110000011101111",
1249=>"00000000000001010000011110010011",
1250=>"11111010111101000010101000100011",
1251=>"00000110100000000000000001101111",
1252=>"11111011110001000010011110000011",
1253=>"00000010000001111000001001100011",
1254=>"11111011010001000010011110000011",
1255=>"00000000000000000000011000010011",
1256=>"11111011110001000010010110000011",
1257=>"00000000000001111000010100010011",
1258=>"11101111100111111110000011101111",
1259=>"00000000000001010000011110010011",
1260=>"11111010111101000010101000100011",
1261=>"00000100000000000000000001101111",
1262=>"00000000000100000000011110010011",
1263=>"11111100111101000010101000100011",
1264=>"00000011010000000000000001101111",
1265=>"11111011110001000010011110000011",
1266=>"00000010000001111000000001100011",
1267=>"11111011010001000010011110000011",
1268=>"11111011010001000000011100010011",
1269=>"00000000000001110000011000010011",
1270=>"11111011110001000010010110000011",
1271=>"00000000000001111000010100010011",
1272=>"11101100000111111110000011101111",
1273=>"00000000110000000000000001101111",
1274=>"00000000000100000000011110010011",
1275=>"11111100111101000010101000100011",
1276=>"00000000000000000000000000010011",
1277=>"11111101010001000010011110000011",
1278=>"00000000000001111001110001100011",
1279=>"11111011010001000010011110000011",
1280=>"11111101000001000010010110000011",
1281=>"00000000000001111000010100010011",
1282=>"10010101100111111111000011101111",
1283=>"00000110110000000000000001101111",
1284=>"11111101000001000010011110000011",
1285=>"00000100010100000000011100010011",
1286=>"00000000111001111010000000100011",
1287=>"11111101000001000010011110000011",
1288=>"00000101001000000000011100010011",
1289=>"00000000111001111010000000100011",
1290=>"11111101000001000010011110000011",
1291=>"00000101001000000000011100010011",
1292=>"00000000111001111010000000100011",
1293=>"11111101000001000010011110000011",
1294=>"00000100111100000000011100010011",
1295=>"00000000111001111010000000100011",
1296=>"11111101000001000010011110000011",
1297=>"00000101001000000000011100010011",
1298=>"00000000111001111010000000100011",
1299=>"00000010110000000000000001101111",
1300=>"11111100000001000010111000100011",
1301=>"11111100110001000010011000000011",
1302=>"11111101000001000010010110000011",
1303=>"11111100100001000010010100000011",
1304=>"11000000000011111111000011101111",
1305=>"11111100110001000010011000000011",
1306=>"11111101000001000010010110000011",
1307=>"11111110110001000010010100000011",
1308=>"11101010000011111111000011101111",
1309=>"00000000000000000000000000010011",
1310=>"00000001100000000000000001101111",
1311=>"11111110000001000010010000100011",
1312=>"10101010100111111111000001101111",
1313=>"00000000000000000000000000010011",
1314=>"10101010000111111111000001101111",
1315=>"00000000000000000000000000010011",
1316=>"10101001100111111111000001101111",

others => (others => '0'));

-- The memory file (use := for an initial value / e.g. program)
shared variable mem : memory_t := prog;

-- Use block RAM for the memory (Xilinx)
attribute ram_style : string;
attribute ram_style of mem : variable is "block";

begin

portA : process (clk)
begin
    if (rising_edge(clk)) then
        dOutA <= mem(to_integer(unsigned(adrA)));
    end if;
end process;

portB : process (clk)
begin
    if (rising_edge(clk)) then

-- Check for write mode
    if (writeEnableB = '1') then
        mem(to_integer(unsigned(adrB))) := dInB;
    end if;
    dOutB <= mem(to_integer(unsigned(adrB)));
-- Synchron read access
    

    end if;
end process;



end Behavioral;